.define res_string_window_title "Startalternativ"
.define res_string_label_ramcard "Kopiera till RAMCard (om det finns)"
.define res_string_label_selector "K|r v{ljare (om s}dan finns)"
