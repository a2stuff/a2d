.define res_string_window_title "Joystick Kalibrering"
.define res_string_label_joy_btn0 "0"
.define res_string_label_joy_btn1 "1"
.define res_string_label_joy_btn2 "2"
