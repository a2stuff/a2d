�~			
	
		



								

	
						                       UU                                                               l68                                                                                                                                                                |                 **                                                               l6l                                                                                                                                                                            UU                                                               8                             66                                                                                                                               < 
     `<<     ** `   X(                 |?||oxoG<?<?>wOoO?<   8               6n                                                                                                                B     ? `BB  6    lUU ` ~~-    0>?3     38ff6ffff0fffff3[fF38f8   0                    ;                                                                                                                  >~  `  ~0l**O0ll l+[   3338033 0y8fff06^CfCffLlL8C8 >>>n6v77;n7>wwwww?                                                                                                              l%  m `
oUUO0~V  +.n -   300<3ml>fs~0v>CfCffLl8xlCl   0f3333n6nn3f3.3fffff3030                                                                                                               ? f%  l?  **gc  6~P[ ?  36333   mlffCf0&vC>C>0fxl80lCl   >f3?3fff3f3f<|<<>3>                                                                                                                %  l ` 
oUUdc   (hs     303033  y|ffCf06fC[f0fx|l0|C|   3f33fff3f3f<|<<333                                                                                                                  ? BB  fl0 l**q~V    +d3   30?033  Fff6fff3ffFfvf3f0F03FfF   3f3333f6ff3f33ff3333                                                                                                               ~   <<  ?l    lUU sll   ~Bn    ?0   |o?<\oo<<O<<0ox?o<o   n;nwoww>>\o?nn                                                                                                                            **        (           0                        0             ?       0       0                                                                                                                                        |?                   UU                                                   `                     3       x                                                                                                                                                               **                                                                                                                                                                                                                                                     UU                                                                                                                                                                                                                                                       **                                                                                                                                                                                                                             