.define res_string_menu_bar_item_file "Arkiv"
.define res_string_menu_bar_item_view "Inneh}ll"
.define res_string_menu_bar_item_special "Speciell"
.define res_string_menu_bar_item_startup "Start"
.define res_string_menu_bar_item_selector "Genv{gar"
.define res_string_menu_item_new_folder "Ny Mapp..."
.define res_char_menu_item_new_folder_shortcut 'N'
.define res_string_menu_item_open "\\ppna"
.define res_char_menu_item_open_shortcut 'O'
.define res_string_menu_item_close "St{ng f|nster"
.define res_char_menu_item_close_shortcut 'W'
.define res_string_menu_item_close_all "St{ng alla"
.define res_string_menu_item_select_all "Markera allt"
.define res_char_menu_item_select_all_shortcut 'A'
.define res_string_menu_item_copy_file "Kopiera en fil..."
.define res_string_menu_item_copy_selection "Kopiera till..."
.define res_string_menu_item_delete_file "Ta bort en fil..."
.define res_string_menu_item_delete_selection "Radera"
.define res_string_menu_item_eject "Mata ut skiva"
.define res_char_menu_item_eject_shortcut 'E'
.define res_string_menu_item_quit "Avsluta"
.define res_char_menu_item_quit_shortcut 'Q'
.define res_string_menu_item_by_icon "Som symboler"
.define res_string_menu_item_by_small_icon "Som sm} symboler"
.define res_string_menu_item_by_name "vid Namn"
.define res_string_menu_item_by_date "efter Datum"
.define res_string_menu_item_by_size "efter Storlek"
.define res_string_menu_item_by_type "efter Typ"
.define res_string_menu_item_check_all_drives "Kontrollera alla enheter"
.define res_string_menu_item_check_drive "Kontrollera Enhet"
.define res_string_menu_item_format_disk "Formatera en disk..."
.define res_string_menu_item_erase_disk "Radera en disk..."
.define res_string_menu_item_disk_copy "Diskkopia..."
.define res_string_menu_item_lock "L}sa..."
.define res_string_menu_item_unlock "L}sa upp..."
.define res_string_menu_item_get_info "Visa info"
.define res_char_menu_item_get_info_shortcut 'I'
.define res_string_menu_item_get_size "F} storlek"
.define res_string_menu_item_rename_icon "Byt namn..."
.define res_string_menu_item_duplicate "Duplicera..."
.define res_string_prompt_button_yes " Ja"
.define res_char_button_yes_shortcut 'J'
.define res_string_prompt_button_no " Nej"
.define res_char_button_no_shortcut 'N'
.define res_string_prompt_button_all " Alla"
.define res_char_button_all_shortcut 'A'
.define res_string_about_text_line5 "F|rfattare: Stephane Cavril, Bernard Gallet, Henri Lamiraux"
.define res_string_about_text_line6 "Richard Danais och Luc Barthelet"
.define res_string_about_text_line7 "Med tack till: A. Gerard, J. Gerber, P. Pahl, J. Bernard"
.define res_string_label_files_remaining "Filer som }terst}r: "
.define res_string_copy_dialog_title "Kopiera..."
.define res_string_copy_label_status "Kopiering: "
.define res_string_copy_label_from "fr}n:"
.define res_string_copy_label_to "till:"
.define res_string_copy_status_files_remaining "Filer som }terst}r att kopiera: "
.define res_string_move_dialog_title "Flytta..."
.define res_string_move_label_status "Flytta: "
.define res_string_move_status_files_remaining "Filer som }terst}r att flytta: "
.define res_string_prompt_overwrite "Den filen finns redan. Vill du skriva |ver det?"
.define res_string_errmsg_too_large_to_copy "Den h{r filen {r f|r stor f|r att kopieras."
.define res_string_errmsg_too_large_to_move "Den h{r filen {r f|r stor f|r att flyttas."
.define res_string_delete_dialog_title "Radera..."
.define res_string_prompt_delete_ok "Klicka p} OK f|r att ta bort: "
.define res_string_label_delete_count "Raderar: "
.define res_string_label_file "Arkiv:"
.define res_string_delete_remaining "Filer som }terst}r att radera: "
.define res_string_delete_prompt_locked_file "Den h{r filen {r l}st, vill du ta bort den {nd}?"
.define res_string_new_folder_label_in "i: "
.define res_string_new_folder_label_name "Nytt mappnamn:"
.define res_string_rename_label_old "Byt namn: "
.define res_string_rename_label_new "Nytt namn:"
.define res_string_rename_label_original "Ursprunglig: "
.define res_string_get_info_label_name "Namn:"
.define res_string_get_info_label_file_size "Storlek:"
.define res_string_get_info_label_create "Skapelsedatum:"
.define res_string_get_info_label_mod "Senaste {ndring:"
.define res_string_get_info_label_type "Typ:"
.define res_string_get_info_label_locked "L}st:"
.define res_string_get_info_label_protected "Skrivskyddad:"
.define res_string_get_info_label_yes "Ja"
.define res_string_get_info_label_no "Nej"
.define res_string_get_info_label_vol_size "Storlek anv{nd/totalt:"
.define res_string_format_disk_label_select "V{lj platsen f|r disken som ska formateras:"
.define res_string_format_disk_label_enter_name "Nytt volymnamn:"
.define res_string_format_disk_prompt_format_prefix "Vill du formatera "
.define res_string_format_disk_prompt_format_suffix "?"
.define res_string_format_disk_status_formatting "Formaterar disken..."
.define res_string_format_disk_error "Formateringsfel. Kontrollera enheten och klicka sedan p} OK f|r att f|rs|ka igen."
.define res_string_erase_disk_label_select "V{lj platsen f|r disken som ska raderas:"
.define res_string_erase_disk_prompt_erase_prefix "Vill du radera "
.define res_string_erase_disk_prompt_erase_suffix "?"
.define res_string_erase_disk_status_erasing "Raderar disken..."
.define res_string_erase_disk_error "Raderingsfel. Kontrollera enheten och klicka sedan p} OK f|r att f|rs|ka igen."
.define res_string_unlock_status_count "Uppl}sning:"
.define res_string_unlock_status_remaining "Filer som }terst}r att l}sa upp: "
.define res_string_lock_status_count "L}sning:"
.define res_string_lock_status_remaining "Filer som }terst}r att l}sa: "
.define res_string_get_size_label_count "Antal filer:"
.define res_string_get_size_label_space "Utrymme som anv{nds p} disk:"
.define res_string_download_dialog_title "Kopiera till RAMCard..."
.define res_string_download_error_ramcard_full "RAMCard {r fullt. Kopian blev inte f{rdig."
.define res_string_warning_insert_system_disk "S{tt i systemdisken."
.define res_string_warning_selector_list_full "Listan {r full. Du m}ste ta bort en genv{g innan du kan l{gga till en ny."
.define res_string_warning_window_must_be_closed "Ett f|nster m}ste st{ngas innan du |ppnar detta f|rem}l."
.define res_string_warning_too_many_files "Det finns f|r m}nga filer f|r att |ppna det h{r objektet!"
.define res_string_warning_too_many_windows "Det finns f|r m}nga f|nster |ppna p} skrivbordet!"
.define res_string_warning_save_changes "Vill du spara {ndringarna p} systemdisken?"
.define res_string_errmsg_00 "Ett ok{nt fel intr{ffade."
.define res_string_errmsg_27 "I/O-fel."
.define res_string_errmsg_28 "Ingen enhet ansluten."
.define res_string_errmsg_2B "Disken {r skrivskyddad."
.define res_string_errmsg_40 "S|kv{gen {r f|r l}ng eller ogiltig."
.define res_string_errmsg_44 "En del av s|kv{gsnamnet finns inte."
.define res_string_errmsg_45 "Volymen kan inte hittas."
.define res_string_errmsg_46 "Filen kan inte hittas."
.define res_string_errmsg_47 "Det namnet finns redan. V{nligen anv{nd ett annat namn."
.define res_string_errmsg_48 "Skivan {r full."
.define res_string_errmsg_49 "Volymkatalogen {r full."
.define res_string_errmsg_4E "Filen {r l}st."
.define res_string_errmsg_52 "Detta {r inte en ProDOS-disk."
.define res_string_errmsg_57 "Det finns en annan volym med det namnet p} skrivbordet."
.define res_string_errmsg_F4 "Att k|ra en bin{r fil kan krascha datorn. [r du s{ker p} att du vill k|ra den?"
.define res_string_errmsg_F5 "En vara kan inte ers{ttas av sig sj{lv eller en vara som den inneh}ller."
.define res_string_errmsg_F6 "Filtyp som inte st|ds."
.define res_string_errmsg_F7 "Det finns inga f|nster |ppna."
.define res_string_errmsg_F8 "Ett objekt kan inte flyttas eller kopieras in i sig sj{lvt."
.define res_string_errmsg_F9 "Det finns 2 volymer med samma namn."
.define res_string_errmsg_FA "Den h{r filen kan inte |ppnas."
.define res_string_errmsg_FB "Det namnet {r f|r l}ngt."
.define res_string_errmsg_FC "V{nligen s{tt i k{lldisken."
.define res_string_errmsg_FD "V{nligen s{tt i destinationsskivan."
.define res_string_errmsg_FE "BASIC.SYSTEM hittades inte."
.define res_string_trash_icon_name "Radera"
.define res_string_sd_prefix_pattern "K#, E#: "
.define res_const_sd_prefix_pattern_offset1 2
.define res_const_sd_prefix_pattern_offset2 6
.define res_string_volume_type_unknown "Ok{nt"
.define res_string_splash_string "Laddar %s..."
.define res_string_prompt_insert_system_disk "S{tt i systemdisken och tryck p} Retur."
.define res_char_resize_shortcut 'G'
.define res_char_move_shortcut 'M'
.define res_char_scroll_shortcut 'X'
.define res_string_auxtype_prefix "     Aux Typ: $"
.define res_string_volume "Volym"
.define res_string_volume_type_disk_ii "Disk II"
.define res_string_volume_type_ramcard "RAMCard"
.define res_string_volume_type_fileshare "AppleShare"
.define res_string_volume_type_vdrive "ADTPro VDRIVE"
.define res_string_selector_label_enter_name "Genv{gsnamn:"
.define res_string_selector_label_add_a_new_entry_to "L{gg till en genv{g till:"
.define res_string_selector_label_primary_run_list "1 meny och lista"
.define res_string_selector_label_secondary_run_list "2 endast lista"
.define res_string_selector_label_download "Kopiera till RAMCard:"
.define res_string_selector_label_at_first_boot "3 vid start"
.define res_string_selector_label_at_first_use "4 vid f|rsta anv{ndningen"
.define res_string_selector_label_never "5 aldrig"
.define res_string_the_dos_33_disk_suffix_pattern "DOS 3.3-skivan i kortplats # enhet #"
.define res_const_the_dos_33_disk_suffix_pattern_offset1 28
.define res_const_the_dos_33_disk_suffix_pattern_offset2 36
.define res_string_the_disk_in_slot_suffix_pattern "disken i kortplats # enhet #"
.define res_const_the_disk_in_slot_suffix_pattern_offset1 20
.define res_const_the_disk_in_slot_suffix_pattern_offset2 28
.define res_string_file_suffix "fil"
.define res_string_files_suffix "filer"
.define res_string_kb_suffix "K"
.define res_string_copy_file_label_source_filename "K{lla filnamn:"
.define res_string_copy_file_label_destination_filename "Destinationsfilnamn:"
.define res_string_delete_file_label_file_to_delete "Fil att radera:"
.define res_string_menu_item_slot_pattern "Kortplats #"
.define res_const_menu_item_slot_pattern_offset1 11
.define res_string_menu_item_add_entry "L{gg till en genv{g..."
.define res_string_menu_item_edit_entry "Redigera en genv{g..."
.define res_string_menu_item_delete_entry "Ta bort en genv{g..."
.define res_string_menu_item_run_entry "K|r en genv{g..."
.define res_string_menu_item_about "Om %s"
.define res_string_window_header_item_suffix " Objekt"
.define res_string_window_header_items_suffix " Objekt"
.define res_string_window_header_k_used_suffix "K i skiva"
.define res_string_window_header_k_available_suffix "K tillg{nglig"
.define res_string_no_date "inget datum"
.define res_string_comma_infix ", "
.define res_string_at_infix " p} "
