�~				
		

						                       UU                                                               66                                                                                                                                                                |                 **                                                               666                                                                                                                                                                            UU                                                                                                                                                                                                                           < 
     `<<     ** `   6    0??     |<??<30cC<<?3CcC?<   0               n                                                                               0                                       B     ? `BB  6    lUU ` >-    33383033     33ff303GGf3f333cccf0f   0                    ;                                                                                8                                        >~  `  0l**O0ll 6k[   300<33 0y3330oOC3C33ss6<C >>3>33333                                                                                                                     l%  6 `
oUUO0~V  .n -   363m63s?0;_C3C33;{6C6   0333333w7333333333030                                                                                                                  ? f%  6?  **gc  6>P; ?  30?033>   m633c30{CC036C6   >33?3333333333>3>                                                                                                                  %  6 ` 
oUUdc   hh     3000330  y>33c30sC03o6>C>   3333333333333333                                                                                                                    ? BB  f60 l**q~V    kd;   3303330  c3ff333cff33gccfc   33333333333333333333                                                                                                                     ~   <<  ?6    lUU sll   >Bn    ?0   |c<?|3c?C<<3cc?c<c   >>>3333>>n3>>>                                                                                                                                         **                                                              ?       0       0       0                                                                                                                                 |?                   UU                                                                                0                                                                                                                                                                **                                                                                                                                                                                                                                                      UU                                                                                                                                                                                                                                                       **                                                                                                                                                                                                                             