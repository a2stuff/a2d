.define res_string_window_title "Ljud"
.define res_string_label_alert "Varningsljud:"
.define res_string_name_silent "Tyst"
.define res_string_name_prodos_buzz "ProDOS Buzz"
.define res_string_name_iigs_bonk "IIgs Bonk"
.define res_string_name_control_g_bell "Control-G Bell"
.define res_string_name_apple_writer_ii "Apple Writer II"
.define res_string_name_dazzle_draw "Dazzle Draw"
.define res_string_name_koala_illustrator "Koala Illustrator"
.define res_string_name_816_paint "816/Paint"
.define res_string_name_apple_panic_1 "Apple Panic 1"
.define res_string_name_apple_panic_2 "Apple Panic 2"
.define res_string_name_bombdrop "Bombdrop"
.define res_string_name_detonate "Detonate"
.define res_string_name_gorgon "Gorgon"
.define res_string_name_versiontel "VersionTel"
.define res_string_name_assembly_line_swoop "Assembly Line Swoop"
.define res_string_name_assembly_line_laser "Assembly Line Laser"
.define res_string_name_assembly_line_bell "Assembly Line Bell"
.define res_string_name_assembly_line_klaxon "Assembly Line Klaxon"
.define res_string_name_obnoxious_whopidoop "Obnoxious Whopidoop"
.define res_string_name_obnoxious_phasor "Obnoxious Phasor"
.define res_string_name_obnoxious_gleep "Obnoxious Gleep"
