.define res_string_window_title "Nyckellayout"
.define res_char_quit_shortcut 'Q'
