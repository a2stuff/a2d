.define res_string_copying_to_ramcard "Kopierar %s till RAMCard..."
.define res_string_label_tip_skip_copying "F|r att hoppa |ver kopiering till RAMCard, h}ll ner \x0F\x1B\x41\x18\x0E n{r du startar."
.define res_string_label_copying "Kopiera till RAMCard: "
.define res_string_prompt_insert_source "S{tt i k{lldisken och tryck p} Retur f|r att forts{tta eller Esc f|r att avbryta."
.define res_string_prompt_ramcard_full "Inte tillr{ckligt med utrymme i RAMCard. Tryck p} Retur f|r att forts{tta."
.define res_string_error_prefix "Fel $"
.define res_string_error_suffix " uppstod vid kopiering "
.define res_string_prompt_copy_not_completed "Kopian blev inte f{rdig. Tryck p} Retur f|r att forts{tta."
.define res_char_monitor_shortcut 'M'
