.define res_filename_calculator Kalkylator
.define res_filename_date_and_time Datum.och.tid
.define res_filename_puzzle Pussel
.define res_filename_sort_directory sortera.katalog
.define res_filename_this_apple detta.apple
.define res_filename_eyes ogon
.define res_filename_screen_dump Skarmdump
.define res_filename_run_basic_here kor.BASIC.har
.define res_filename_key_caps nyckellayout
.define res_filename_find_files hitta.filer
.define res_filename_control_panels kontrollpaneler
.define res_filename_control_panel kontrollpanel
.define res_filename_options alternativ
.define res_filename_system_speed systemhastighet
.define res_filename_joystick styrspak
.define res_filename_international Internationellt
.define res_filename_screen_savers skarmslackare
.define res_filename_toys Leksaker
.define res_filename_flying_toasters brodrostar
.define res_filename_neko Neko
.define res_filename_map Karta
.define res_filename_melt smalta
.define res_filename_matrix matrix
.define res_filename_invert negativ
.define res_filename_calendar Kalender
.define res_filename_sounds Ljud
.define res_filename_analog_clock analog.klocka
.define res_filename_digital_clock digital.klocka
.define res_filename_print_catalog Skriv.katalog
