 	 > |     >>  <    U*               ??3?>333?3333?33   0               33  A?  @ AA  B   	 *U ?@    0   333333?33333333330   0                     @ @ ]]wU*`66  ?    !3333?7333333333 ># * @ >@$EUR
 0 w*UN1I        -?3;?3;3333333   033++030  @kk@&EM>
? ! U*?d?!        =333333333303??3?   >33++>3> * @? >@?]U
 0 w*Uq?!   ?	      3333333333333?3333   333++333   @AA  
 U*{~j           3?3?3?33333?33   ?>+?? *   |  @>>  O     *U  66                             >                0                                             0         z     U*                                                                                              