.define res_string_window_title "Alternativ"
.define res_string_label_ramcard "Kopiera till RAMCard (om det finns)"
.define res_string_label_selector "K|r Selector vid start"
.define res_string_label_shortcuts "Visa genv{gar i dialogrutor"
