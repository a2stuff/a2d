.define res_string_button_fixed "Fast teckenbredd"
.define res_string_button_prop "Proportionerligt"
