.define res_string_window_title "Ljud"
.define res_string_label_alert "Varningsljud:"
.define res_string_name_silent "Tyst"
