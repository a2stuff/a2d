.define res_string_dc_menu_bar_item_file "Arkiv"
.define res_string_menu_bar_item_facilities "Alternativ"
.define res_string_dc_menu_item_quit "Avsluta"
.define res_char_dc_menu_item_quit_shortcut 'Q'
.define res_string_menu_item_quick_copy "Snabb Kopia"
.define res_string_dc_menu_item_disk_copy "Diskkopia"
.define res_string_button_read_drive "L{s Drives"
.define res_char_button_read_drive_shortcut 'D'
.define res_string_label_slot_drive_name "Kortplats, Enhet, Namn"
.define res_string_prompt_select_source "V{lj k{lldisk"
.define res_string_prompt_select_destination "V{lj destinationsskiva"
.define res_string_label_status_formatting "Formaterar disken..."
.define res_string_label_status_writing "Skrivande...   "
.define res_string_label_status_reading "L{sning...    "
.define res_string_unknown "Ok{nt"
.define res_string_label_select_quit "V{lj Avsluta fr}n Arkiv-menyn (%cQ) f|r att g} tillbaka till skrivbordet"
.define res_string_label_blocks_read "Block L{s: "
.define res_string_label_blocks_written "Block skrivna: "
.define res_string_label_blocks_to_transfer "Block att |verf|ra: "
.define res_string_source "K{lla "
.define res_string_destination "Destination "
.define res_string_slot_prefix "Kortplats "
.define res_string_drive_infix "  Diskenhet "
.define res_string_dos33_s_d_pattern "DOS 3.3 K#, E# "
.define res_const_dos33_s_d_pattern_offset1 10
.define res_const_dos33_s_d_pattern_offset2 14
.define res_string_dos33_disk_copy "DOS 3.3 diskkopia"
.define res_string_pascal_disk_copy "Pascal skiva kopia"
.define res_string_prodos_disk_copy "ProDOS diskkopia"
.define res_string_escape_stop_copy " Esc stoppa kopian"
.define res_string_error_writing "Fel vid skrivblock "
.define res_string_error_reading "Fel vid l{sning av block "
.define res_string_prompt_insert_source "S{tt i k{lldisken och klicka p} OK."
.define res_string_prompt_insert_destination "S{tt i m}lskivan och klicka p} OK."
.define res_string_prompt_erase_prefix "Vill du radera "
.define res_string_prompt_erase_suffix "?"
.define res_string_errmsg_dest_format_fail "M}lskivan kan inte formateras!"
.define res_string_errmsg_format_error "Fel under formatering."
.define res_string_errmsg_dest_protected "Destinationsvolymen {r skrivskyddad!"
.define res_string_prompt_erase_slot_drive_pattern "Vill du radera disken i kortplats # enhet #?"
.define res_const_prompt_erase_slot_drive_pattern_offset1 35
.define res_const_prompt_erase_slot_drive_pattern_offset2 43
.define res_string_label_status_copy_success "Kopian lyckades."
.define res_string_label_status_copy_fail "Kopian blev inte f{rdig."
.define res_string_prompt_insert_source_or_cancel "S{tt i k{llskivan eller tryck p} Esc f|r att avbryta."
.define res_string_prompt_insert_dest_or_cancel "S{tt i m}lskivan eller tryck p} Esc f|r att avbryta."
