.define res_string_label_find "S|k:"
.define res_string_button_search "S|k          \x0D"
