�~							
                       UU                                                                                                                                                                                                                                  |                 **                                                                                                                                                                                                                                            UU                                                                                              
                                                                                                                                < 
      <<     ** _    
         <A!!A!A                  

&                                                                                                                            B       BB     	 UU _  %	         B"	"	c#""!A!""
                                                                                                                                                     >~      	**oll 
	   
   9U%AA!"A 	%A                                                                                                                             $%  
 @
wUUo~  
F    	%1I%AA!"A   [A
                                                                                                                           ? "%  
  **wA  
)      %"!A)AA!"A"   I
*                                                                                                                           ?%  
 @ 
wUUv	A   *       y>!A)A]!*>A>   I
*                                                                                                                                BB  "
  **y~    ))         A"	"	A1""	!D!A"A   	I
                                                                                                                            ~   <<  
    UU {ll   F       <A<A!\D!AA   I                                                                                                                                                **                                                              ?                                                                                                                                                       |?                   UU                                                                                                                                                                                                                                                    **                                                                                                                                                                                                                                                       UU                                                                                                                                                                                                                                                        **                                                                                                                                                                                                                              