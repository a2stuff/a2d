.define res_filename_calculator "Kalkylator"
.define res_filename_date_and_time "Datum.och.Tid"
.define res_filename_puzzle "Pussel"
.define res_filename_lights_out "Lights.Out"
.define res_filename_sort_directory "Sortera.Katalog"
.define res_filename_eyes "Ogon"
.define res_filename_print_screen "Utskrift.Skarm"
.define res_filename_screenshot "Skarmdump"
.define res_filename_run_basic_here "Kor.BASIC.Har"
.define res_filename_key_caps "Nyckellayout"
.define res_filename_find_files "Hitta.Filer"
.define res_filename_control_panels "Kontrollpaneler"
.define res_filename_control_panel "Kontrollpanel"
.define res_filename_options "Alternativ"
.define res_filename_system_speed "Systemhastighet"
.define res_filename_joystick "Styrspak"
.define res_filename_international "Internationellt"
.define res_filename_screen_savers "Skarmslackare"
.define res_filename_toys "Leksaker"
.define res_filename_flying_toasters "Brodrostar"
.define res_filename_helix "Helix"
.define res_filename_bounce "Studsa"
.define res_filename_neko "Neko"
.define res_filename_map "Karta"
.define res_filename_melt "Smalta"
.define res_filename_matrix "Matrix"
.define res_filename_invert "Negativ"
.define res_filename_random "Slumpmassigt"
.define res_filename_rods_pattern "Rods.Pattern"
.define res_filename_calendar "Kalender"
.define res_filename_sounds "Ljud"
.define res_filename_analog_clock "Analog.Klocka"
.define res_filename_digital_clock "Digital.Klocka"
.define res_filename_print_catalog "Skriv.Katalog"
.define res_filename_change_type "Andra.Typ"
.define res_filename_benchmark "Benchmark"
.define res_filename_message "Meddelande"
.define res_filename_cd_remote "CD.Fjarr"
.define res_filename_darkness "Morker"
.define res_filename_round_corners "Runda.Horn"
.define res_filename_sci_calc "Sci.Berakn"
.define res_filename_dos33_import "DOS33.Importera"
.define res_filename_views "Innehallen"
.define res_filename_this_apple "This.Apple"
.define res_filename_show_text_file "Show.Text.File"
.define res_filename_show_image_file "Show.Image.File"
.define res_filename_show_duet_file "Show.Duet.File"
.define res_filename_show_font_file "Show.Font.File"
