.define res_string_error_string "Fel "
.define res_string_window_title "Kalkylator"
