.define res_string_window_title "Studsa"
