.define res_string_message_placeholder "Skriv ett meddelande..."
