.define res_string_select_disk "Select DOS 3.3 disk:"
.define res_string_slot_drive_pattern "Slot #  Drive #"
.define res_const_slot_drive_pattern_offset1 6
.define res_const_slot_drive_pattern_offset2 15
.define res_string_disk_volume_prefix "Disk Volume "
.define res_string_button_import "Importera"
