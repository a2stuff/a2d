.define res_string_select_disk "V{lj DOS 3.3-disk:"
.define res_string_slot_drive_pattern "Kortplats #  Diskenhet #"
.define res_const_slot_drive_pattern_offset1 11
.define res_const_slot_drive_pattern_offset2 24
.define res_string_disk_volume_prefix "Disk Volume "
.define res_string_button_import "Importera"
