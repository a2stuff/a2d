.define res_string_window_title "Alternativ"
.define res_string_label_ramcard "Kopiera till RAMCard (om det finns)"
.define res_string_label_selector "Visa Genv{gar vid start"
.define res_string_label_shortcuts "Visa kortkommandon i dialogrutor"
.define res_string_label_case "Bevara versaler och gemener i namn"
.define res_string_label_invisible "Visa osynliga filer"
