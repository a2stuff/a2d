�~				
		
		
	



		
                       UU                                                               ll8                                                                                                                                                                |                 **                                                               lll                               8                                                                                                                                             UU                                                               8                             l6l                                                                                                                               < 
     `<<     ** `   6X     0<0>     |x:z<:1nn::FnNxx   0               l68n                                                                                                                 B     ? `BB  ,   lUU ` 6~K    0666066     ll&LFl5<jY,ll,}YY2l,l   0 <                   ;                                                                            8                                      >~  `  0l**O0ll 6l.-   6063 yfl#L&nX4X<X~l0l4Xp1f~f <<4<[;<67768<<                                                                                                                  l-  6 `
oUUO0~V  
+    63m6<LfL6llLf606LLL0L6f6   6666666mm6666mm=6d666                                                                                                             ? f-  6?  **gc  6h} ?  ?0   m3fFf|<lL38LlL0L333   333336ll>66ll623>3                                                                                                                  -  6 ` 
oUUdc   4g     0  y;ffclf6f36lfff8f0;3;   36636666:3                                                                                                                       ? BB  &60 l**q~V    R3     {3c3ff6f3fv6vlV{{   66366a                                                                                                                    ~   <<  6   lUU sll   `N       <N_|?|^F~Fv6Fvc;LFl|NN   vv>v~?~qq3cwv8^vlv~|vv                                                                                                                        **                                                       P    ?                    6                                                                                                                               |?                   UU                                                          `                                                                                                                                                                                 **                                                                                                                                                                                                                                                      UU                                                                                                                                                                                                                                                       **                                                                                                                                                                                                                             