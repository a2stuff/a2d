.define res_string_label_date_separator "Datumavgr{nsare:"
.define res_string_label_time_separator "Tidsavgr{nsare:"
.define res_string_label_decimal_separator "Decimalavgr{nsare:"
.define res_string_label_thousands_separator "Tusentalsavgr{nsare:"
