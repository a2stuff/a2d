�~				
			

						                       UU                                                               33                                                                                                                                                                |                 **                                                               33                                                                                                                                                                            UU                                                                                            33                                                                                                                               < 
     `     ** `   6    ???3?????     ????????303_??????33Cc3????   0 <              33_                                                                                                                     B     ? `      lUU ` [-    3003033     036630[[333333Cc30333?   0                    [                                                                                                                       >~  `==  0l**O0ll 6?   3003033< 0}36630[[333333C6303333 ???????????????33C33????{                                                                                                                      l%  6 `
oUUO0~V   -   3?????0??<m?>6;?0[[3?3??33C???3?  033333[333333C30030                                                                                                                    ? f=  6?  **gc  6s ?  30003030   <m366330C[33033[333   ?33?33[3333?3[3??3?                                                                                                                     =  6 ` 
oUUdc   h|c     30003030  }366333C[33033[6333   33333[333303[3333                                                                                                                       ?   60 l**q~V    hZs   30003030<  366333C[3303[c333   33333[333303[3333                                                                                                                  ~     ?6    lUU sll   x    ???0??0??   3?????3?3?C{??3??c?3?3   ??????33[3????<?3?????                                                                                                                                      **                                                             ?       0       0       0                                                                                                                                 |?                   UU                                                                        ?       0       ?                                                                                                                                                         **                                                                                                                                                                                                                                                      UU                                                                                                                                                                                                                                                       **                                                                                                                                                                                                                             