.define res_string_window_title "Inst{llningspanelen"
.define res_string_label_pattern "Skrivbordsm|nster"
.define res_string_label_rgb_color "RGB-f{rg"
.define res_string_label_dblclick_speed "Dubbelklicka p} Speed"
.define res_string_label_mouse_tracking "Mussp}rning"
.define res_string_label_slow "L}ngsam"
.define res_string_label_fast "Snabb"
.define res_string_label_ipblink1 "Ins{ttningspunkten"
.define res_string_label_ipblink2 "blinkar"
