.define res_string_button_ok "OK"
.define res_string_button_cancel "Avbryt"
.define res_string_button_cancel_shortcut "Esc"
.define res_string_button_try_again "F|rs|k igen"
.define res_char_button_try_again_shortcut 'F'
.define res_string_button_yes "Ja"
.define res_char_button_yes_shortcut 'J'
.define res_string_button_no "Nej"
.define res_char_button_no_shortcut 'N'
.define res_string_button_all "Alla"
.define res_char_button_all_shortcut 'A'
.define res_string_shortcut_apple_1 " (\x1F1)"
.define res_string_shortcut_apple_2 " (\x1F2)"
.define res_string_shortcut_apple_3 " (\x1F3)"
.define res_string_shortcut_apple_4 " (\x1F4)"
.define res_string_shortcut_apple_5 " (\x1F5)"
.define res_string_shortcut_apple_6 " (\x1F6)"
.define res_char_shortcut_resize 'G'
.define res_char_shortcut_move 'M'
.define res_char_shortcut_scroll 'X'
.define res_char_shortcut_close 'W'
.define res_string_button_drives "Enheter"
.define res_string_button_open "\\ppna"
.define res_string_button_close "St{ng"
.define res_string_shortcut_drives "^D"
.define res_string_shortcut_open "^O"
.define res_string_shortcut_close "^C"
.define res_string_copyright_line1 "Copyright Apple Computer Inc., 1986"
.define res_string_copyright_line2 "Copyright Version Soft, 1985 - 1986"
.define res_string_copyright_line3 "Alla r{ttigheter f|rbeh}lls"
.define res_string_prompt_insert_system_disk "S{tt i systemdisken och tryck p} Retur."
.define res_string_weekday_abbrev_1 "Sol"
.define res_string_weekday_abbrev_2 "M}n"
.define res_string_weekday_abbrev_3 "Tis"
.define res_string_weekday_abbrev_4 "Ons"
.define res_string_weekday_abbrev_5 "Tor"
.define res_string_weekday_abbrev_6 "Fre"
.define res_string_weekday_abbrev_7 "L|r"
.define res_string_month_name_1 "Januari"
.define res_string_month_name_2 "Februari"
.define res_string_month_name_3 "Mars"
.define res_string_month_name_4 "April"
.define res_string_month_name_5 "Maj"
.define res_string_month_name_6 "Juni"
.define res_string_month_name_7 "Juli"
.define res_string_month_name_8 "Augusti"
.define res_string_month_name_9 "September"
.define res_string_month_name_10 "Oktober"
.define res_string_month_name_11 "November"
.define res_string_month_name_12 "December"
.define res_string_month_abbrev_1 "Jan"
.define res_string_month_abbrev_2 "Feb"
.define res_string_month_abbrev_3 "Mar"
.define res_string_month_abbrev_4 "Apr"
.define res_string_month_abbrev_5 "Maj"
.define res_string_month_abbrev_6 "Jun"
.define res_string_month_abbrev_7 "Jul"
.define res_string_month_abbrev_8 "Aug"
.define res_string_month_abbrev_9 "Sep"
.define res_string_month_abbrev_10 "Okt"
.define res_string_month_abbrev_11 "Nov"
.define res_string_month_abbrev_12 "Dec"
.define res_char_decimal_separator ','
.define res_char_thousands_separator ' '
.define res_char_date_separator '-'
.define res_char_time_separator '.'
.define res_const_date_order 1
.define res_const_clock_format 128
.define res_string_version_format_long "%s Version %d.%d%s"
.define res_string_noprod_version_format_long "Version %d.%d%s"
