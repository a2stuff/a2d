          ?  ?           
 ?                                                                                                  <                 
** ?                                                                                                 ?    
 /          33                  .  " >  6 
**/ 7      3                           6 
7            ? 6?  **7   ?                
:              >     
**9    ;          ??           
 ;

          33
   3
     <                
** ?                                                                                                               
 ?                                                                                                    ?  ?            ** ?                                                                                                   