.define res_string_window_title "\\gon"
