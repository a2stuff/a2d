.define res_string_window_title "Om denna Apple II"
.define res_string_model_ii "Apple ]["
.define res_string_model_iiplus "Apple ][+"
.define res_string_model_iii "Apple /// (efterliknande)"
.define res_string_model_iie_original "Apple IIe (ursprunglig)"
.define res_string_model_iie_enhanced "Apple IIe F|rb{ttras"
.define res_string_model_iie_edm "Apple IIe (EDM)"
.define res_string_model_iie_card "Apple IIe Option Card"
.define res_string_model_iic_original "Apple //c (ROM 255)"
.define res_string_model_iic_rom0 "Apple //c (ROM 0)"
.define res_string_model_iic_rom3 "Apple //c (ROM 3)"
.define res_string_model_iic_rom4 "Apple //c (ROM 4)"
.define res_string_model_iic_plus "Apple IIc Plus"
.define res_string_model_iigs_pattern "Apple IIgs (ROM #)"
.define res_const_model_iigs_pattern_offset1 17
.define res_string_model_laser128 "Laser 128"
.define res_string_model_ace500 "Franklin ACE 500"
.define res_string_model_ace2000 "Franklin ACE 2X00"
.define res_string_model_tlc "Tiger Learning Computer"
.define res_string_model_trackstar_e "Trackstar E"
.define res_string_model_trackstar_plus "Trackstar Plus"
.define res_string_model_mega_iie "Mega IIe"
.define res_string_model_tk3000 "Microdigital TK-3000 //e"
.define res_string_model_pravetz "Pravetz 8A/C"
.define res_string_prodos_version_pattern "ProDOS #.#.#"
.define res_const_prodos_version_pattern_offset1 8
.define res_const_prodos_version_pattern_offset2 10
.define res_const_prodos_version_pattern_offset3 12
.define res_string_slot_n_pattern "Kortplats #:   "
.define res_const_slot_n_pattern_offset1 11
.define res_string_memory_prefix "Minne: "
.define res_string_memory_kb_suffix "K"
.define res_string_memory_mb_suffix "MB"
.define res_string_card_type_diskii "Disk II"
.define res_string_card_type_block "Generic Block Device"
.define res_string_card_type_smartport "SmartPort: "
.define res_string_card_type_ssc "Super Serial Card"
.define res_string_card_type_80col "80 Kolumn Kort"
.define res_string_card_type_mouse "Muskort"
.define res_string_card_type_silentype "Silentype"
.define res_string_card_type_clock "Klocka"
.define res_string_card_type_comm "Kommunikationskort"
.define res_string_card_type_serial "Seriekort"
.define res_string_card_type_parallel "Parallellt Kort"
.define res_string_card_type_printer "Skrivarkort"
.define res_string_card_type_joystick "Styrspak"
.define res_string_card_type_io "I/O-Kort"
.define res_string_card_type_modem "Modem"
.define res_string_card_type_audio "Ljudkort"
.define res_string_card_type_storage "Masslagring"
.define res_string_card_type_network "N{tverkskort"
.define res_string_card_type_mockingboard "Mockingboard"
.define res_string_card_type_z80 "Z-80 Kort"
.define res_string_card_type_uthernet2 "Uthernet II"
.define res_string_card_type_lcmeve "Le Chat Mauve Eve"
.define res_string_card_type_vidhd "VidHD"
.define res_string_card_type_grappler "Grappler Parallel Printer Card"
.define res_string_card_type_thunderclock "ThunderClock"
.define res_string_card_type_applecat "Apple-CAT II Modem"
.define res_string_card_type_workstation "Workstation Card"
.define res_string_device_type_cricket "The Cricket!"
.define res_string_device_type_nvram "NVRAM Block Device"
.define res_string_device_type_booti "BOOTI Block Device"
.define res_string_unknown "(ok{nt)"
.define res_string_empty "(t|mma)"
.define res_string_none "(ingen)"
.define res_string_duplicate_suffix_pattern " (#)"
.define res_const_duplicate_suffix_pattern_offset1 3
.define res_string_cpu_prefix "    CPU: "
.define res_string_cpu_type_6502 "6502"
.define res_string_cpu_type_65C02 "65C02"
.define res_string_cpu_type_65C02zip "65C02 (ZIP CHIP)"
.define res_string_cpu_type_R65C02 "R65C02"
.define res_string_cpu_type_65802 "65802"
.define res_string_cpu_type_65816 "65816"
.define res_char_easter_egg_shortcut 'E'
