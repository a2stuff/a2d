.define res_string_label_clock_12hour "12 tim"
.define res_string_label_clock_24hour "24 tim"
