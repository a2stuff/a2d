 	 > ?w     >>  <    U*   68      8??     ??3?<333?33333?33   0               33   A?!  @ AA  B    *U ?@ 63   `333<3033   6!333330?333333333330   0 &                       @ ]]w>U*`66 ?0   0;006330-3330?73333333336 >>>6>;>33#33>>> *   >@$EUR 0 w*UN1I   0> > ?30> =3;?03;33333   37#3337+3373'33+30333&  kk@&EM>? ! U*?d?!  [ 0   70?033   333330333303?333   333?33+333333+3333*  ? >@?]U 0 w*Uq?!   ?33  3303333  ?3333333333333?3?3?   ;3#;;3+333;0&;+;3;  ?- @AA   U*{~j  0n 8   ??0   >3?>3?3?33333?33   76>63<6<+3663>77 *   ?  @>>  O     *U  66                                              0                    0       0                 w0         z     U*                                                                                0             