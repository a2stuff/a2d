.define res_string_window_title "CPU Benchmark (MHz)"
.define res_string_60hz "60Hz"
.define res_string_50hz "50Hz"
