.define res_string_status_loading_desktop "Startar Apple II DeskTop..."
.define res_string_menu_bar_item_file "Arkiv"
.define res_string_menu_bar_item_edit "Redigera"
.define res_string_menu_bar_item_view "Inneh}ll"
.define res_string_menu_bar_item_special "Speciell"
.define res_string_menu_bar_item_startup "Start"
.define res_string_menu_bar_item_selector "Genv{gar"
.define res_string_menu_item_new_folder "Ny Mapp"
.define res_char_menu_item_new_folder_shortcut 'N'
.define res_string_menu_item_open "\\ppna"
.define res_char_menu_item_open_shortcut 'O'
.define res_string_menu_item_close "St{ng"
.define res_string_menu_item_close_all "St{ng alla"
.define res_string_menu_item_select_all "Markera allt"
.define res_char_menu_item_select_all_shortcut 'A'
.define res_string_menu_item_copy_selection "Kopiera till..."
.define res_string_menu_item_delete_selection "Radera"
.define res_string_menu_item_eject "Mata ut skiva"
.define res_char_menu_item_eject_shortcut 'E'
.define res_string_menu_item_quit "Avsluta"
.define res_char_menu_item_quit_shortcut 'Q'
.define res_string_menu_item_cut "Klipp ut"
.define res_char_menu_item_cut_shortcut 'X'
.define res_string_menu_item_copy "Kopiera"
.define res_char_menu_item_copy_shortcut 'C'
.define res_string_menu_item_paste "Klistra in"
.define res_char_menu_item_paste_shortcut 'V'
.define res_string_menu_item_clear "Rensa"
.define res_string_menu_item_by_icon "Som symboler"
.define res_string_menu_item_by_small_icon "Som sm} symboler"
.define res_string_menu_item_by_name "vid Namn"
.define res_string_menu_item_by_date "efter Datum"
.define res_string_menu_item_by_size "efter Storlek"
.define res_string_menu_item_by_type "efter Typ"
.define res_string_menu_item_check_all_drives "Kontrollera alla enheter"
.define res_string_menu_item_check_drive "Kontrollera Enhet"
.define res_string_menu_item_format_disk "Formatera disk..."
.define res_string_menu_item_erase_disk "Radera disk..."
.define res_string_menu_item_disk_copy "Kopia disk ..."
.define res_string_menu_item_make_link "Skapa alias"
.define res_string_menu_item_show_original "Visa original"
.define res_string_menu_item_get_info "Visa info"
.define res_char_menu_item_get_info_shortcut 'I'
.define res_string_menu_item_rename_icon "Byt namn"
.define res_string_menu_item_duplicate "Duplicera"
.define res_char_menu_item_duplicate_shortcut 'D'
.define res_string_new_folder_default "New.Folder"
.define res_string_about_text_line5 "F|rfattare: Stephane Cavril, Bernard Gallet, Henri Lamiraux"
.define res_string_about_text_line6 "Richard Danais och Luc Barthelet"
.define res_string_about_text_line7 "Med tack till: A. Gerard, J. Gerber, P. Pahl, J. Bernard"
.define res_string_label_files_remaining "Filer som }terst}r: "
.define res_string_copy_label_status "Kopiering: "
.define res_string_copy_label_from "fr}n:"
.define res_string_copy_label_to "till:"
.define res_string_move_label_status "Flytta: "
.define res_string_prompt_overwrite "Den filen finns redan. Vill du byta ut den?"
.define res_string_error_unknown "Ett ok{nt fel intr{ffade."
.define res_string_error_too_large_to_copy "Den h{r filen {r f|r stor f|r att kopieras."
.define res_string_error_too_large_to_move "Den h{r filen {r f|r stor f|r att flyttas."
.define res_string_error_overwrite_dir "En mapp kan inte ers{ttas av ett annat objekt. Radera det sedan f|rs|k igen."
.define res_string_prompt_delete_confirm_singular_format "[r du s{ker p} att du vill ta bort %0n fil permanent?"
.define res_string_prompt_delete_confirm_plural_format "[r du s{ker p} att du vill ta bort %0n filer permanent?"
.define res_string_label_delete_count "Raderar: "
.define res_string_label_file "Arkiv:"
.define res_string_delete_prompt_locked_file "Den h{r filen {r l}st, vill du ta bort den {nd}?"
.define res_string_get_info_label_name "Namn:"
.define res_string_get_info_label_file_size "Storlek:"
.define res_string_get_info_label_create "Skapad:"
.define res_string_get_info_label_mod "[ndrad:"
.define res_string_get_info_label_type "Typ:"
.define res_string_get_info_checkbox_locked "L}st"
.define res_string_get_info_shortcut_locked " (^L)"
.define res_string_get_info_label_protected "Skrivskyddad:"
.define res_string_get_info_label_yes "Ja"
.define res_string_get_info_label_no "Nej"
.define res_string_get_info_label_vol_size "Storlek anv{nd/totalt:"
.define res_string_get_info_size_file_format "%0k"
.define res_string_get_info_size_dir_singular_format "%0k f|r %1n objekt  "
.define res_string_get_info_size_dir_plural_format "%0k f|r %1n objekt  "
.define res_string_get_info_size_vol_singular_format "%0k f|r %1n objekt / %2k  "
.define res_string_get_info_size_vol_plural_format "%0k f|r %1n objekt / %2k  "
.define res_string_format_disk_label_select "V{lj platsen f|r disken som ska formateras:"
.define res_string_format_disk_label_location "Platsen: "
.define res_string_format_disk_label_enter_name "Nytt volymnamn:"
.define res_string_format_disk_status_formatting "Formaterar disken..."
.define res_string_format_disk_error "Formateringsfel. Kontrollera enheten."
.define res_string_erase_disk_label_select "V{lj platsen f|r disken som ska raderas:"
.define res_string_erase_disk_prompt_erase_format "[r du s{ker att du vill radera %0s?"
.define res_string_erase_disk_status_erasing "Raderar disken..."
.define res_string_erase_disk_error "Raderingsfel. Kontrollera enheten."
.define res_string_tip_copy_prodos "Tips: Kopiera PRODOS till disken f|r att g|ra den startbar."
.define res_string_download_error_ramcard_full "RAMCard {r fullt. Kopian blev inte f{rdig."
.define res_string_alert_selector_list_full "Listan {r full. Du m}ste ta bort en genv{g innan du kan l{gga till en ny."
.define res_string_alert_window_must_be_closed "Ett f|nster m}ste st{ngas innan du |ppnar detta f|rem}l."
.define res_string_alert_too_many_files "Det finns f|r m}nga filer f|r att |ppna det h{r objektet!"
.define res_string_alert_too_many_windows "Det finns f|r m}nga f|nster |ppna p} skrivbordet!"
.define res_string_alert_save_changes "Vill du spara {ndringarna p} systemdisken?"
.define res_string_alert_confirm_running "Att k|ra en bin{r fil kan krascha datorn. [r du s{ker p} att du vill k|ra den?"
.define res_string_alert_bad_replacement "En vara kan inte ers{ttas av sig sj{lv eller en vara som den inneh}ller."
.define res_string_alert_unsupported_type "Filtyp som inte st|ds."
.define res_string_alert_no_windows_open "Det finns inga f|nster |ppna."
.define res_string_alert_move_copy_into_self "Ett objekt kan inte flyttas eller kopieras in i sig sj{lvt."
.define res_string_alert_duplicate_volume_names "Det finns 2 volymer med samma namn."
.define res_string_alert_cannot_open "Den h{r filen kan inte |ppnas."
.define res_string_alert_name_too_long "Det namnet {r f|r l}ngt."
.define res_string_alert_unreadable_format "Den h{r disken kunde inte l{sas. Vill du formatera det?"
.define res_string_trash_icon_name "Radera"
.define res_string_sd_name_format "K%0d, E%1d: %2s"
.define res_string_volume_type_unknown "Ok{nt"
.define res_string_auxtype_format "%0s         Aux Typ: $%1x"
.define res_string_folder "Mapp"
.define res_string_volume "Volym"
.define res_string_volume_type_disk_ii "Disk II"
.define res_string_volume_type_ramcard "RAMCard"
.define res_string_volume_type_fileshare "AppleShare"
.define res_string_volume_type_vdrive "ADTPro VDRIVE"
.define res_string_selector_label_enter_name "Genv{gsnamn:"
.define res_string_selector_label_add_a_new_entry_to "Visa genv{g i:"
.define res_string_selector_label_primary_run_list "meny och lista"
.define res_string_selector_label_secondary_run_list "endast lista"
.define res_string_selector_label_download "Kopiera till RAMCard:"
.define res_string_selector_label_at_first_boot "vid start"
.define res_string_selector_label_at_first_use "vid f|rsta anv{ndningen"
.define res_string_selector_label_never "aldrig"
.define res_string_the_dos_33_disk_format "DOS 3.3-skivan i kortplats %0d enhet %1d"
.define res_string_the_disk_in_slot_format "disken i kortplats %0d enhet %1d"
.define res_string_file_count_singular_format "%0n fil"
.define res_string_file_count_plural_format "%0n filer"
.define res_string_kb_suffix "K"
.define res_string_menu_item_slot_pattern "Kortplats #"
.define res_const_menu_item_slot_pattern_offset1 11
.define res_string_menu_item_add_entry "L{gg till en genv{g..."
.define res_string_menu_item_edit_entry "Redigera en genv{g..."
.define res_string_menu_item_delete_entry "Ta bort en genv{g..."
.define res_string_menu_item_run_entry "K|r en genv{g..."
.define res_string_menu_item_about "Om Apple II DeskTop"
.define res_string_menu_item_about_this_apple "Om denna Apple II"
.define res_string_window_header_item_count_singular_format "%0n Objekt"
.define res_string_window_header_item_count_plural_format "%0n Objekt"
.define res_string_window_header_k_used_format "%0k i skiva"
.define res_string_window_header_k_available_format "%0k tillg{nglig"
.define res_string_no_date "inget datum"
.define res_string_datetime_format "%0s p} %1s"
.define res_string_mdy_format "%1s %0d, %2d"
.define res_string_dmy_format "%0d %1s %2d"
.define res_string_today "Idag"
.define res_string_yesterday "Ig}r"
.define res_string_tomorrow "Imorgon"
