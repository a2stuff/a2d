.define res_string_playing "Spelar: "
.define res_string_credit1 "Electric Duet av Paul Lutus"
.define res_string_credit2 "Musikspelare av Alexander Patalenski och Cybernesto"
.define res_string_instructions "Tryck p} valfri tangent f|r att avbryta"
