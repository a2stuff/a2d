.define res_string_button_norm "Normal          N"
.define res_char_button_norm_shortcut 'N'
.define res_string_button_fast "Snabb          S"
.define res_char_button_fast_shortcut 'S'
.define res_string_dialog_title "Systemhastighet"
