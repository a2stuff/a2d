.define res_string_label_type "Typ:  $"
.define res_string_label_auxtype "Aux Typ:  $"
.define res_string_err_no_files_selected "Det finns inga filer valda."
