.define res_string_label_type "Typ:  $"
.define res_string_label_auxtype "Aux Typ:  $"
