.define res_string_selector_name "Genv{gar"
.define res_string_status_loading_selector "Startar Genv{gar..."
.define res_string_alert_selector_unable_to_run "Det g}r inte att k|ra programmet."
.define res_string_alert_io_error "I/O-fel."
.define res_string_alert_no_device "Ingen enhet ansluten."
.define res_string_alert_pathname_does_not_exist "En del av s|kv{gsnamnet finns inte."
.define res_string_alert_insert_source_disk "V{nligen s{tt i k{lldisken."
.define res_string_alert_file_not_found "Filen kan inte hittas."
.define res_string_alert_insert_system_disk "S{tt i systemdisken."
.define res_string_alert_basic_system_not_found "BASIC.SYSTEM hittades inte."
.define res_string_menu_bar_item_file "Arkiv"
.define res_string_menu_bar_item_startup "Start"
.define res_string_menu_item_run_a_program "K|r ett program..."
.define res_char_menu_item_run_a_program_shortcut 'R'
.define res_string_menu_item_slot_pattern "Kortplats #"
.define res_const_menu_item_slot_pattern_offset1 11
.define res_string_button_desktop "Skrivbord"
.define res_char_button_desktop_shortcut 'S'
.define res_string_label_download "Kopierar till RAMCard..."
.define res_string_label_copying "Kopierar: "
.define res_string_errmsg_not_enough_room "Inte tillr{ckligt med utrymme i RAMCard f|r att kopiera programmet."
.define res_string_errmsg_copy_incomplete "Ett fel uppstod under nedladdningen. Kopian blev inte f{rdig."
.define res_string_label_files_to_copy "Filer att kopiera: "
.define res_string_label_files_remaining "Filer som }terst}r: "
